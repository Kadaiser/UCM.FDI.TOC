`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:06:51 10/21/2015 
// Design Name: 
// Module Name:    rec_patron_baba 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module rec_patron_baba(
    input entrada STD_LOGIC;
    output salida STD_LOGIC
    );


endmodule
